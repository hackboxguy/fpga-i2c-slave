`define VERSION_MAGIC_START 16'hAE25
`define VERSION_MAGIC_END   16'hE025
`define VERSION_MAJOR       8'd1
`define VERSION_MINOR       8'd0
`define BUILD_NUMBER        16'd42
`define GIT_COMMIT_HASH_HI  16'hDEAD
`define GIT_COMMIT_HASH_LO  16'hBEEF
`define BUILD_TIMESTAMP_HI  16'h690E
`define BUILD_TIMESTAMP_LO  16'h5186
`define I2C_SLAVE_ADDRESS   7'h3A
`define VERSION_BRAM_SIZE   16
`define VERSION_BRAM_DEPTH  8
